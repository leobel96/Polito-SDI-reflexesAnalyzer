LIBRARY ieee;
USE ieee.std_logic_1164.all; 

ENTITY voter IS 
	PORT
	(
		Q_RX_REG :  IN  STD_LOGIC_VECTOR (7 DOWNTO 0);
		VOTER_OUT :  OUT STD_LOGIC
	);
END ENTITY voter;

ARCHITECTURE structural OF voter IS 
BEGIN
	VOTER_OUT <= (Q_RX_REG(4) AND Q_RX_REG(5) AND Q_RX_REG(6)) OR (Q_RX_REG(3) AND Q_RX_REG(5) AND Q_RX_REG(6)) OR 
					 (Q_RX_REG(3) AND Q_RX_REG(4) AND Q_RX_REG(6)) OR (Q_RX_REG(3) AND Q_RX_REG(4) AND Q_RX_REG(5)) OR 
					 (Q_RX_REG(2) AND Q_RX_REG(5) AND Q_RX_REG(6)) OR (Q_RX_REG(2) AND Q_RX_REG(4) AND Q_RX_REG(6)) OR
					 (Q_RX_REG(2) AND Q_RX_REG(4) AND Q_RX_REG(5)) OR (Q_RX_REG(2) AND Q_RX_REG(3) AND Q_RX_REG(6)) OR 
					 (Q_RX_REG(2) AND Q_RX_REG(3) AND Q_RX_REG(5)) OR (Q_RX_REG(2) AND Q_RX_REG(3) AND Q_RX_REG(4));					 
END ARCHITECTURE structural;
